entity CSAdder is
  port (
    
  ) ;
end CSAdder;

architecture arch of CSAdder is



begin



end architecture ; -- arch