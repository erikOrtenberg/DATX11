entity MUX is
  port (
    
  ) ;
end MUX ;

architecture arch of MUX is



begin



end architecture ; -- arch